ROMBLOCK_inst : ROMBLOCK PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
